`ifndef TEST_OVERRIDE_DEFS_VH
`define TEST_OVERRIDE_DEFS_VH

`define RX_PAYLOAD_Q_SIZE_W 3
`define RX_PAYLOAD_Q_SIZE   (2**`RX_PAYLOAD_Q_SIZE_W)
`define PAYLOAD_BUF_MEM_ELS (`MAX_FLOW_CNT * `RX_PAYLOAD_Q_SIZE)
`define PAYLOAD_BUF_MEM_ADDR_W (`BSG_SAFE_CLOG2(`PAYLOAD_BUF_MEM_ELS))
`define PAYLOAD_ENTRY_ADDR_W 16
`define PAYLOAD_ENTRY_LEN_W 8

`define MAX_FLOW_CNT 8
`endif