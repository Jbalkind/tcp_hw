`ifndef SIM_CONFIG
`define SIM_CONFIG

`define REAL_REMOTE
//`define CYCLE_LOG
`endif
