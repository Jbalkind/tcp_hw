`ifndef TEST_OVERRIDE_DEFS_VH
`define TEST_OVERRIDE_DEFS_VH

`define     MAX_FLOW_CNT            8// should be power of two

`define     PAYLOAD_ENTRY_ADDR_W 16
`define     PAYLOAD_ENTRY_LEN_W 8

`define PAYLOAD_PTR_W  16
`define RX_PAYLOAD_PTR_W `PAYLOAD_PTR_W
`endif
